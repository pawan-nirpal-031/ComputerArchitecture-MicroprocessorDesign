module full_adder(sum,cout,a,b,cin);
    output sum,cout;
    input a,b,cin;
    wire x,y,z;
    

endmodule